// Module Name: mips_single_cycle_datapath.v
// Project: MIPS Single Cycle Processor
// Description: Datapath module.
// Author: Cengiz Mert ÖNCE
// Date: 2026-01-09

module mips_single_cycle_datapath
(
    input wire clk,
    input wire reset,
    input wire [31:0] instruction, // Instruction provided as input
    output wire [31:0] alu_result, // ALU output
    output wire [31:0] write_data  // Data written to register
);

wire [5:0] opcode;      // instruction[31:26]
wire [4:0] rs;          // instruction[25:21]
wire [4:0] rt;          // instruction[20:16]
wire [4:0] rd;          // instruction[15:11]
wire [4:0] shamt;       // instruction[10:6] (not used)
wire [5:0] funct;       // instruction[5:0]
wire [15:0] immediate;  // instruction[15:0]
    
// Map instruction fields to named wires
assign opcode    = instruction[31:26];
assign rs        = instruction[25:21];
assign rt        = instruction[20:16];
assign rd        = instruction[15:11];
assign shamt     = instruction[10:6];
assign funct     = instruction[5:0];
assign immediate = instruction[15:0];

// ----------------
// Control Signals wires
wire RegDst;        // Selects between rt and rd for write register
wire Branch;        // Branch control signal
wire MemRead;      // Memory read control signal
wire MemtoReg;     // Selects between ALU result and memory data for write data
wire [1:0] ALUOp;       // ALU operation control signal
wire MemWrite;    // Memory write control signal
wire ALUSrc;       // Selects between register data and immediate for ALU input
wire RegWrite;     // Register write control signal

// Control Unit instance
control_unit CU (
    .opcode(opcode),
    .reg_dst(RegDst),
    .alu_src(ALUSrc),
    .reg_write(RegWrite),
    .alu_op(ALUOp)
);
// ----------------

// Register File wires
wire [31:0] read_data1; // Data from register rs
wire [31:0] read_data2; // Data from register rt
wire [4:0] write_register; // Data from rs or rt based on instruction type 

mux2to1_5bit rt_rd_write_reg_mux (
    .in0(rt),          // I-type instruction uses rt
    .in1(rd),          // R-type instruction uses rd
    .sel(RegDst),      // Control signal to select between rt and rd
    .y(write_register)  // Output write register
);


// register file instance
register_file RF (
    .clk(clk),
    .reset(reset),
    .reg_write(RegWrite),
    .read_reg1(rs),
    .read_reg2(rt),
    .write_reg(write_register[4:0]),
    .write_data(write_data),

    .read_data1(read_data1),
    .read_data2(read_data2)
);

// Sign Extender instance
// ALU input 2 selection
wire [31:0] extended_immediate;

sign_extender SE (
    .immediate_in(immediate),
    .immediate_out(extended_immediate)
);

wire [31:0] alu_input2;
para_mux2to1 #(.DATA_WIDTH(32)) ALU_second_src_mux (
    .inputA(read_data2),            // Register data (rt)
    .inputB(extended_immediate),    // Sign-extended immediate
    .select(ALUSrc),                // Control signal to select ALU input
    .outputY(alu_input2)                      // ALU input 2
);

// ALU control signal generation
wire [3:0] alu_control_out; // ALU control signal - generated by ALU control unit
alu_control ALU_CTRL (
    .alu_op(ALUOp),
    .funct(funct),
    .alu_control(alu_control_out) // ALU control signal
);

// ALU instance
wire alu_zero;
alu ALU (
    .a(read_data1),                 // ALU input 1 (from register rs)
    .b(alu_input2),                 // ALU input 2 (from mux)
    .alu_control(alu_control_out),  // ALU control signal
    .result(alu_result),            // ALU result output
    .zero(alu_zero)                 // Zero flag (not used here)
);

// assign write_data = alu_result; // if we wanna write alu result to register

endmodule